const string _NULL_STRING = "";
const byte   _DOT = ".";
