`ifndef _NULL_STRING
`define _NULL_STRING
const string _NULL_STRING = "";
`endif

`ifndef _DOT
`define _DOT
const byte   _DOT = ".";
`endif
