const string _NULL_STRING = "";
