`ifndef __MOCK_UVM_COMPARER__
`define __MOCK_UVM_COMPARER__

import uvm_pkg::*;

class mock_uvm_comparer extends uvm_comparer;
endclass

`endif
