import uvm_pkg::*;

class uvm_boat_anchor;
endclass
